= next require './next'
:= (require './numbers') a b

console.log (next a)
console.log (next b)
