= numbers | 1 2 3

|= numbers first second third

console.log first
console.log second
console.log third
