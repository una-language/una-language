= add
  -> first
    -> second
      + first second

= addOne add 1

>> (addOne 3)
