= numbers | 1 2 3

|= numbers first second third

>> first
>> second
>> third
