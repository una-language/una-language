console.log true
console.log false

console.log (! true)
console.log (! false)

console.log (&& true true true)
console.log (&& true false true)
console.log (|| false false false)
console.log (|| false true false)
