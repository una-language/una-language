= a (+ 1 2 3)
= b +
  1
  2
  3
= c + 1
  2
  3

console.log a
console.log b
console.log c
