= x 1
= greeting "Hello World!"
