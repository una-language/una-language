= object :
  a 1
  b :
    c 2
    d 3
  e 4
  f 5

:= object a (b c d) e f

>_ a
>_ c
>_ d
>_ e
>_ f
