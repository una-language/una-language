console.log
  ? true 1 0

console.log
  ? (> 2 1) 'Greater' 'Less'

console.log
  ? (> 2 1)
    ? (> 1 2) 'x' 'y'
    'z'
