--> './constant'
--> './string'
--> './array'
--> './object'
--> './function'
--> './module'
