= numbers | 1 2 3

|= numbers first second third

>_ first
>_ second
>_ third
