= add
  -> first
    -> second
      + first second

= addOne add 1

>_ (addOne 3)
