console.log '--------------------- Constant ---------------------'

= number 1
console.log number
