= next (--> './next')
:= (--> './numbers') a b

>_ (next a)
>_ (next b)
