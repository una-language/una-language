= integer 4

>_ integer
>_ (- integer)
>_ (+ integer 1)
>_ (- integer 1)
>_ (* integer 2)
>_ (/ integer 2)
>_ (% integer 3)

= float 4.5

>_ float
>_ (- float)
>_ (+ float 1.2)
>_ (- float 1.2)
>_ (* float 3)
>_ (/ float 1.5)
