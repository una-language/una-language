= next -> number
  + number 1

module.exports next
