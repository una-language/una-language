= users |
  :
    name 'Alice'
    age 20
  : (name 'Bob') (age 25)


console.log users
console.log (.0 users)
