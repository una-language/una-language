--> 1
