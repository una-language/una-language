= digits | 0 1 2 3 4 5 6 7 8 9

>> digits

>>
  | 1 2 3

= numbers |
  12
  34
  57
  93

>> numbers

>>
  numbers.get 0

>>
  numbers.length

>>
  numbers.size

= numbersWithFirstElementAdded numbers.addFirst 0
= numbersWithLastElementAdded numbers.addLast 123
= numbersWithElementAdded numbers.add 145

>> numbersWithFirstElementAdded
>> numbersWithLastElementAdded
>> numbersWithElementAdded
