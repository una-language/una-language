console.log 'Constant declaration'
console.log '-----------'
=-> './constant-declaration'
console.log '-----------\n'

console.log 'Numbers'
console.log '-----------'
=-> './numbers'
console.log '-----------\n'

console.log 'Comparison'
console.log '-----------'
=-> './comparison'
console.log '-----------\n'

console.log 'Condition'
console.log '-----------'
=-> './condition'
console.log '-----------\n'

console.log 'Function'
console.log '-----------'
=-> './function'
console.log '-----------\n'

console.log 'List'
console.log '-----------'
=-> './list'
console.log '-----------\n'

console.log 'Map'
console.log '-----------'
=-> './map'
console.log '-----------\n'

console.log 'Average age'
console.log '-----------'
=-> './average-age'
console.log '-----------\n'
