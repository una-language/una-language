= integer 4

console.log integer
console.log - integer
console.log + integer 1
console.log - integer 1
console.log * integer 2
console.log / integer 2
console.log % integer 3

= float 4.5

console.log float
console.log - float
console.log + float 1.2
console.log - float 1.2
console.log * float 3
console.log / float 1.5


console.log + 1 2 3
console.log - 8 2 1
console.log * 3 4 5
console.log / 16 2 2
