= name 'John'

console.log
 'Hello ${name}!'
