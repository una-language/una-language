= pet
  -> (voice food)
    :
      voice
      food

= cat pet 'Meow' 'Milk'
= dog pet 'Woof' 'Meat'

>_ cat
>_ dog
