console.log
  + 2 2

console.log
  - 6 2

console.log
  * 2 2

console.log
  / 8 2

console.log
  / 10 2.5
