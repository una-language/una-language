= digits | 0 1 2 3 4 5 6 7 8 9

console.log digits

|= digits zero one two
console.log zero
console.log one
console.log two

= numbers |
  12
  34
  57
  93

console.log numbers

console.log (numbers.get 0)

console.log (numbers.size)

console.log (numbers.addFirst 0)
console.log (numbers.addLast 123)
console.log (numbers.add 145)
