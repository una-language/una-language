console.log
  ? true 1 0

console.log
  ? (> 2 1) 'ok' 'not ok'

console.log
  ? (> 2 1)
    ? (> 1 2) 'x' 'y'
    'z'
