console.log '--------------------- Module ---------------------'

= data --> './data'

console.log data.first
console.log (data.addSecond 4)
