= integer 4

console.log integer
console.log (- integer)
console.log (+ integer 1)
console.log (- integer 1)
console.log (* integer 2)
console.log (/ integer 2)
console.log (% integer 3)

= float 4.5

console.log float
console.log (- float)
console.log (+ float 1.2)
console.log (- float 1.2)
console.log (* float 3)
console.log (/ float 1.5)
