>_ 'Single quoted string with "text inside double quotes"'
>_ "Double quoted string with 'text inside single quotes'"

= planet 'Earth'
>_ 'Hello ${planet}!'

= text `
  'First line of text'
  'Second line of text'
  'Third line of text'

>_ text
