= a :
  b :
    c 1

>_
  ?. a.b.c

>_
  ?. a.b.d

>_
  ?. a.d.e
