console.log
  ' (Hello World!)
