<-- 1
