--> './next' next
--> './numbers' numbers

:= numbers a b

console.log (next a)
console.log (next b)
