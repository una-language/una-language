= next -> number (+ number 1)

<- next
