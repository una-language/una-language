>_ 'Hello'
>_ "Hello World!"

= string 'Hello World!'
>_ string

= name 'John'
= greeting 'Hello ${name}'
>_ greeting

= text `
  'First line of text'
  'Second line of text'
  'Third line of text'

>_ text
