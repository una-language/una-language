= x >= 2 3

console.log x
