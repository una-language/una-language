>_ (> 2 1)
>_ (< 1 2)
>_ (>= 1 1)
>_ (<= 1 1)
>_ (== 1 "1")
>_ (=== 1 1)
>_ (!= 1 2)
>_ (!== 1 "1")

>_
  ? (> 2 1) 15 30
