= number <-
  = three (+ 1 2)
  * three 4

console.log number
