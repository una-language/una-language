>> 'Hello World!'
