<-- :
  first (--> './first')
  addSecond -> (. number) (+ number (--> './second'))
