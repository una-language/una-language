= object :
  b :
    c 2.0

console.log object.b
