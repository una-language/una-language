= e 3

= object :
  a 1
  b :
    c 2.0
    d 'Hello'
  e
  f | 4 5 6

>_ object
>_ object.a
>_ object.b
>_ object.b.c
>_ object.b.d
>_ object.e
>_ object.f
