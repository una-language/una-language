=-> './data' (: greeting name)
=-> './handler' handle

handle greeting name
