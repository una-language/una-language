= a <- 'a'
= b 'b'

console.log a
console.log b
