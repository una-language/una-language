= integer 4

>> integer
>> (- integer)
>> (+ integer 1)
>> (- integer 1)
>> (* integer 2)
>> (/ integer 2)
>> (% integer 3)

= float 4.5

>> float
>> (- float)
>> (+ float 1.2)
>> (- float 1.2)
>> (* float 3)
>> (/ float 1.5)


>> (+ 1 2 3)
>> (- 8 2 1)
>> (* 3 4 5)
>> (/ 16 2 2)
