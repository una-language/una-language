= object :
  a 1
  b :
    c 2
    d 3
  e 4
  f 5

= numbers | 1 2 3

console.log numbers
