= first true
= second false

>_ first
>_ second
>_
  ! second

>_
  && true true true

>_
  && true false true

>_
  || false false false

>_
  || false true false
