= greeting 'Hello World!'

>> greeting
