>> 'Single quoted string with "text inside double quotes"'
>> "Double quoted string with 'text inside single quotes'"

= planet 'Earth'
>> 'Hello ${planet}!'

= text `
  'First line of text'
  'Second line of text'
  'Third line of text'

>> text
