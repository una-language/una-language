= digits | 0 1 2 3 4 5 6 7 8 9

>> digits

|= digits zero one two
>> zero
>> one
>> two

= numbers |
  12
  34
  57
  93

>> numbers

>> numbers.get 0

>> numbers.length
>> numbers.size

>> numbers.addFirst 0
>> numbers.addLast 123
>> numbers.add 145
