= sum
  -> (first second)
    + first second

console.log (sum 1 2)
