= object :
  a 1
  b :
    c 2

= (: a ( b : c:d )) object
console.log a
console.log d
