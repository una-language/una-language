= a 1

= b --
  = one 1
  + one 1

= c <-
  = oneAndHalf 1.5
  * oneAndHalf 2

= d -> number
  = eight 8
  / eight number

>> a
>> b
>> c
>> (d 2)
