= digits | 0 1 2 3 4 5 6 7 8 9

console.log digits

console.log
  | 1 2 3

= numbers |
  12
  34
  57
  93

console.log numbers

console.log
  numbers.get 0

console.log
  numbers.length

console.log
  numbers.size

= numbersWithFirstElementAdded numbers.addFirst 0
= numbersWithLastElementAdded numbers.addLast 123
= numbersWithElementAdded numbers.add 145

console.log numbersWithFirstElementAdded
console.log numbersWithLastElementAdded
console.log numbersWithElementAdded
