console.log 'Average age'
console.log '-----------'
=-> './average-age'
console.log '-----------'
