>> 'Hello'
>> "Hello World!"

= string 'Hello World!'
>> string

= name 'John'
= greeting 'Hello ${name}'
>> greeting

= text `
  'First line of text'
  'Second line of text'
  'Third line of text'

>> text
