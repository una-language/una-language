console.log '--------------------- Array ---------------------'

= numbers . 1 2 3 4
console.log numbers

= (. first second ...rest) numbers
console.log first
console.log second
console.log rest
