= greeting 'Hello World!'

>_ greeting
