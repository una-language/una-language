>> (> 2 1)
>> (< 1 2)
>> (>= 1 1)
>> (<= 1 1)
>> (== 1 "1")
>> (=== 1 1)
>> (!= 1 2)
>> (!== 1 "1")

>>
  ? (> 2 1) 15 30
