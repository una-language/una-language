= object :
  a 1
  b :
    c 2.0
    d 'Hello'
  e 3
  f | 4 5 6

console.log object
console.log object.a
console.log object.b
console.log object.b.c
console.log object.b.d
console.log object.e
console.log object.f
