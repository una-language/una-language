console.log
  ' (Hello world!)
