= add
  -> first
    -> second
      + first second

= addOne add 1

console.log
  addOne 3
