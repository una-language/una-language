= numbers | 1 2 3

console.log numbers
