= next (--> './next')
:= (--> './numbers') a b

>> (next a)
>> (next b)
