console.log 'Hello World!'
