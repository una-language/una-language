= numbers | 1 2 3 4

= result
  numbers.map
    -> number :
      a number
      b number

console.log result
