= list | 1 2 3 4

console.log list
console.log
  list.map (-> x (+ x 1))

= (| first second) list

console.log first
console.log second
