require './constant'
require './array'
require './object'
require './function'
