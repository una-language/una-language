= a :
  b :
    c 1

>>
  ?. a.b.c

>>
  ?. a.b.d

>>
  ?. a.d.e
