<-- 2
