<-= -> (greeting name)
  console.log greeting
  console.log name
