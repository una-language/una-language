>_ 'Hello World!'
