--> './next' next

console.log (next 2)
