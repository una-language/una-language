--> 2
