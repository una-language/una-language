<-- './constant'
<-- './string'
<-- './array'
<-- './object'
<-- './function'
<-- './module'
<-- './fizzbuzz'
