= first true
= second false

>> first
>> second
>>
  ! second

>>
  && true true true

>>
  && true false true

>>
  || false false false

>>
  || false true false
