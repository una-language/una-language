= object :
  b :
    c 2.0

>> object.b
