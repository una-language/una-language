console.log 'Constant declaration'
console.log '-----------'
=-> './constant-declaration'
console.log '-----------\n'

console.log 'Numbers'
console.log '-----------'
=-> './numbers'
console.log '-----------\n'

console.log 'Comparison'
console.log '-----------'
=-> './comparison'
console.log '-----------\n'

console.log 'Average age'
console.log '-----------'
=-> './average-age'
console.log '-----------\n'
