= object :
  a 1
  b :
    c 2
    d 3
  e 4
  f 5

:= object a (b c d) e f

console.log a
console.log c
console.log d
console.log e
console.log f
