= x ? (> 2 1) (<- null)

console.log x
