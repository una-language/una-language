= a :
  b 'g'

console.log a
console.log a.b
console.log (a.b.toString ())
