= digits | 0 1 2 3 4 5 6 7 8 9

>_ digits

>_
  | 1 2 3

= numbers |
  12
  34
  57
  93

>_ numbers

>_
  numbers.get 0

>_
  numbers.length

>_
  numbers.size

= numbersWithFirstElementAdded numbers.addFirst 0
= numbersWithLastElementAdded numbers.addLast 123
= numbersWithElementAdded numbers.add 145

>_ numbersWithFirstElementAdded
>_ numbersWithLastElementAdded
>_ numbersWithElementAdded
