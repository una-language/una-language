= x (+ 1 2)

console.log x
