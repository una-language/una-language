= first --> './first'
= second --> './second'

<-- :
  first
  addSecond -> (. number) (+ number second)
