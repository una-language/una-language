console.log (> 2 1)
console.log (< 1 2)
console.log (>= 1 1)
console.log (<= 1 1)
console.log (== 1 "1")
console.log (=== 1 1)
console.log (!= 1 2)
console.log (!== 1 "1")

console.log
  ? (> 2 1) 15 30
