= number 1
console.log number
